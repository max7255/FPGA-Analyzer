`timescale 	100ps / 100ps
//-------------------------------------
// GAMMA_8_12.v
//-------------------------------------
// History of Changes:
//	6-16-2009  Initial creation
//-------------------------------------
// This module applies a fixed gamma to a video path
//-------------------------------------
// Programmed with a gamma of 2.2
// Latency is 1 cycle.
//-------------------------------------
module GAMMA_8_12 (
input	wire			CLK,  // Master Clock
input	wire			CE,   // clock enable
input	wire			EN,   // if no enable, a gamma of 1.0 is applied.
input	wire	[7:0]	DIN,
output	wire	[11:0]	DOUT
);

wire	[15:0]	gamma_out;
assign DOUT = gamma_out[11:0];
RAMB16_S18 #(
	// Address 0 to 255 are gamma 1.0 for no EN
	.INIT_00(256'h00f0_00e0_00d0_00c0_00b0_00a0_0090_0080_0070_0060_0050_0040_0030_0020_0010_0000),
	.INIT_01(256'h01f1_01e1_01d1_01c1_01b1_01a1_0191_0181_0171_0161_0151_0141_0131_0121_0111_0101),
	.INIT_02(256'h02f2_02e2_02d2_02c2_02b2_02a2_0292_0282_0272_0262_0252_0242_0232_0222_0212_0202),
	.INIT_03(256'h03f3_03e3_03d3_03c3_03b3_03a3_0393_0383_0373_0363_0353_0343_0333_0323_0313_0303),
	.INIT_04(256'h04f4_04e4_04d4_04c4_04b4_04a4_0494_0484_0474_0464_0454_0444_0434_0424_0414_0404),
	.INIT_05(256'h05f5_05e5_05d5_05c5_05b5_05a5_0595_0585_0575_0565_0555_0545_0535_0525_0515_0505),
	.INIT_06(256'h06f6_06e6_06d6_06c6_06b6_06a6_0696_0686_0676_0666_0656_0646_0636_0626_0616_0606),
	.INIT_07(256'h07f7_07e7_07d7_07c7_07b7_07a7_0797_0787_0777_0767_0757_0747_0737_0727_0717_0707),
	.INIT_08(256'h08f8_08e8_08d8_08c8_08b8_08a8_0898_0888_0878_0868_0858_0848_0838_0828_0818_0808),
	.INIT_09(256'h09f9_09e9_09d9_09c9_09b9_09a9_0999_0989_0979_0969_0959_0949_0939_0929_0919_0909),
	.INIT_0A(256'h0afa_0aea_0ada_0aca_0aba_0aaa_0a9a_0a8a_0a7a_0a6a_0a5a_0a4a_0a3a_0a2a_0a1a_0a0a),
	.INIT_0B(256'h0bfb_0beb_0bdb_0bcb_0bbb_0bab_0b9b_0b8b_0b7b_0b6b_0b5b_0b4b_0b3b_0b2b_0b1b_0b0b),
	.INIT_0C(256'h0cfc_0cec_0cdc_0ccc_0cbc_0cac_0c9c_0c8c_0c7c_0c6c_0c5c_0c4c_0c3c_0c2c_0c1c_0c0c),
	.INIT_0D(256'h0dfd_0ded_0ddd_0dcd_0dbd_0dad_0d9d_0d8d_0d7d_0d6d_0d5d_0d4d_0d3d_0d2d_0d1d_0d0d),
	.INIT_0E(256'h0efe_0eee_0ede_0ece_0ebe_0eae_0e9e_0e8e_0e7e_0e6e_0e5e_0e4e_0e3e_0e2e_0e1e_0e0e),
	.INIT_0F(256'h0fff_0fef_0fdf_0fcf_0fbf_0faf_0f9f_0f8f_0f7f_0f6f_0f5f_0f4f_0f3f_0f2f_0f1f_0f0f),
	// Address 256 to 511 are gamma 2.2
	.INIT_10(256'h0008_0007_0006_0005_0004_0003_0003_0002_0002_0001_0001_0000_0000_0000_0000_0000), 
	.INIT_11(256'h0028_0025_0022_0020_001D_001B_0019_0017_0015_0013_0011_000F_000E_000C_000B_0009), 
	.INIT_12(256'h0063_005F_005A_0056_0052_004D_0049_0046_0042_003E_003B_0037_0034_0031_002E_002B), 
	.INIT_13(256'h00BD_00B6_00B0_00AA_00A4_009E_0098_0092_008C_0087_0081_007C_0077_0072_006D_0068), 
	.INIT_14(256'h0137_012E_0126_011E_0115_010D_0105_00FE_00F6_00EE_00E7_00E0_00D8_00D1_00CA_00C4), 
	.INIT_15(256'h01D3_01C8_01BD_01B3_01A8_019E_0194_018A_0180_0177_016D_0164_015B_0151_0148_0140), 
	.INIT_16(256'h0291_0284_0277_026B_025E_0252_0245_0239_022D_0221_0216_020A_01FF_01F4_01E8_01DD), 
	.INIT_17(256'h0374_0364_0355_0346_0337_0329_031A_030C_02FE_02F0_02E2_02D4_02C6_02B9_02AB_029E), 
	.INIT_18(256'h047B_046A_0458_0447_0436_0425_0414_0403_03F3_03E2_03D2_03C2_03B2_03A2_0392_0383), 
	.INIT_19(256'h05A9_0595_0581_056D_055A_0546_0533_0520_050D_04FA_04E8_04D5_04C3_04B1_049F_048D), 
	.INIT_1A(256'h06FD_06E6_06D0_06BA_06A4_068E_0679_0663_064E_0639_0624_060F_05FA_05E5_05D1_05BD), 
	.INIT_1B(256'h0878_085F_0847_082E_0816_07FD_07E5_07CD_07B6_079E_0786_076F_0758_0741_072A_0713), 
	.INIT_1C(256'h0A1C_0A01_09E6_09CA_09AF_0995_097A_0960_0945_092B_0911_08F7_08DE_08C4_08AB_0891), 
	.INIT_1D(256'h0BE9_0BCB_0BAD_0B8F_0B72_0B54_0B37_0B1A_0AFD_0AE1_0AC4_0AA8_0A8C_0A6F_0A54_0A38), 
	.INIT_1E(256'h0DDF_0DBE_0D9E_0D7E_0D5D_0D3E_0D1E_0CFE_0CDF_0CBF_0CA0_0C81_0C62_0C44_0C25_0C07), 
	.INIT_1F(256'h0FFF_0FDC_0FB9_0F96_0F73_0F50_0F2E_0F0C_0EEA_0EC8_0EA6_0E84_0E63_0E42_0E21_0E00)
	) gammalut (
	.CLK(CLK),    // Clock
	.ADDR({1'b0, EN, DIN[7:0]}),  // 10-bit Address Input
	.DO(gamma_out), .DOP(), 
	.DI(16'h0000), .DIP(2'b00), .WE(1'b0), 
	.EN(CE), .SSR(1'b0)
	);

endmodule
