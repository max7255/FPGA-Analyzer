`timescale 	100ps / 100ps
//-------------------------------------
// INV_GAMMA_12_8.v
//-------------------------------------
// History of Changes:
//	6-16-2009  Initial creation
//-------------------------------------
// This module applies a fixed inverse gamma to a video path
//-------------------------------------
// Programmed with a gamma of 1/2.2
// Latency is 2 cycles.
//-------------------------------------
module INV_GAMMA_12_8 (
input	wire			CLK,  // Master Clock
input	wire			CE,   // clock enable
input	wire			EN,   // if no enable, a gamma of 1.0 is applied.
input	wire	[11:0]	DIN,
output	reg 	[7:0]	DOUT
);

// Implemented with two 8-bit wide RAMB16's - High and Low
// It would have been technically better to have used 2 4-wide parts, 
// which would span the full 4k address space, 
// but the INIT's would not have been as clear, and we have a mux stage
// on the output anyway for the !EN bypass mode, so no big performance 
// or resource hit here.
wire	[7:0]	gamma_outL, gamma_outH;
// Lower half of table
RAMB16_S9 #(
	// Address 0 to 511
	.INIT_00(256'h1C_1B_1B_1A_1A_1A_19_19_18_18_17_17_16_16_15_15_14_13_13_12_11_11_10_0F_0E_0D_0C_0B_0A_08_06_00), 
	.INIT_01(256'h26_26_26_25_25_25_25_24_24_24_23_23_23_22_22_22_21_21_21_20_20_20_1F_1F_1F_1E_1E_1E_1D_1D_1C_1C), 
	.INIT_02(256'h2E_2E_2E_2D_2D_2D_2D_2D_2C_2C_2C_2C_2B_2B_2B_2B_2A_2A_2A_2A_29_29_29_29_28_28_28_28_27_27_27_27), 
	.INIT_03(256'h35_34_34_34_34_34_33_33_33_33_33_32_32_32_32_32_31_31_31_31_31_30_30_30_30_30_2F_2F_2F_2F_2F_2E), 
	.INIT_04(256'h3A_3A_3A_3A_3A_39_39_39_39_39_39_38_38_38_38_38_38_37_37_37_37_37_36_36_36_36_36_36_35_35_35_35), 
	.INIT_05(256'h3F_3F_3F_3F_3F_3F_3E_3E_3E_3E_3E_3E_3D_3D_3D_3D_3D_3D_3D_3C_3C_3C_3C_3C_3C_3B_3B_3B_3B_3B_3B_3A), 
	.INIT_06(256'h44_44_44_44_43_43_43_43_43_43_43_42_42_42_42_42_42_42_41_41_41_41_41_41_40_40_40_40_40_40_40_3F), 
	.INIT_07(256'h48_48_48_48_48_48_47_47_47_47_47_47_47_46_46_46_46_46_46_46_46_45_45_45_45_45_45_45_44_44_44_44), 
	.INIT_08(256'h4C_4C_4C_4C_4C_4C_4B_4B_4B_4B_4B_4B_4B_4B_4A_4A_4A_4A_4A_4A_4A_4A_49_49_49_49_49_49_49_49_48_48), 
	.INIT_09(256'h50_50_50_50_4F_4F_4F_4F_4F_4F_4F_4F_4F_4E_4E_4E_4E_4E_4E_4E_4E_4D_4D_4D_4D_4D_4D_4D_4D_4D_4C_4C), 
	.INIT_0A(256'h53_53_53_53_53_53_53_53_53_52_52_52_52_52_52_52_52_52_52_51_51_51_51_51_51_51_51_50_50_50_50_50), 
	.INIT_0B(256'h57_57_57_57_56_56_56_56_56_56_56_56_56_56_55_55_55_55_55_55_55_55_55_54_54_54_54_54_54_54_54_54), 
	.INIT_0C(256'h5A_5A_5A_5A_5A_5A_59_59_59_59_59_59_59_59_59_59_58_58_58_58_58_58_58_58_58_58_57_57_57_57_57_57), 
	.INIT_0D(256'h5D_5D_5D_5D_5D_5D_5D_5D_5C_5C_5C_5C_5C_5C_5C_5C_5C_5C_5B_5B_5B_5B_5B_5B_5B_5B_5B_5B_5A_5A_5A_5A), 
	.INIT_0E(256'h60_60_60_60_60_60_60_60_5F_5F_5F_5F_5F_5F_5F_5F_5F_5F_5E_5E_5E_5E_5E_5E_5E_5E_5E_5E_5E_5D_5D_5D), 
	.INIT_0F(256'h63_63_63_63_63_63_62_62_62_62_62_62_62_62_62_62_62_62_61_61_61_61_61_61_61_61_61_61_61_60_60_60), 
	// Address 512 to 1023
	.INIT_10(256'h66_66_66_66_65_65_65_65_65_65_65_65_65_65_65_65_64_64_64_64_64_64_64_64_64_64_64_63_63_63_63_63), 
	.INIT_11(256'h68_68_68_68_68_68_68_68_68_68_68_68_67_67_67_67_67_67_67_67_67_67_67_67_66_66_66_66_66_66_66_66), 
	.INIT_12(256'h6B_6B_6B_6B_6B_6B_6B_6B_6A_6A_6A_6A_6A_6A_6A_6A_6A_6A_6A_6A_69_69_69_69_69_69_69_69_69_69_69_69), 
	.INIT_13(256'h6E_6E_6D_6D_6D_6D_6D_6D_6D_6D_6D_6D_6D_6D_6D_6C_6C_6C_6C_6C_6C_6C_6C_6C_6C_6C_6C_6B_6B_6B_6B_6B), 
	.INIT_14(256'h70_70_70_70_70_70_70_70_6F_6F_6F_6F_6F_6F_6F_6F_6F_6F_6F_6F_6F_6E_6E_6E_6E_6E_6E_6E_6E_6E_6E_6E), 
	.INIT_15(256'h72_72_72_72_72_72_72_72_72_72_72_72_72_71_71_71_71_71_71_71_71_71_71_71_71_71_71_70_70_70_70_70), 
	.INIT_16(256'h75_75_75_75_75_74_74_74_74_74_74_74_74_74_74_74_74_74_73_73_73_73_73_73_73_73_73_73_73_73_73_73), 
	.INIT_17(256'h77_77_77_77_77_77_77_77_77_76_76_76_76_76_76_76_76_76_76_76_76_76_76_75_75_75_75_75_75_75_75_75), 
	.INIT_18(256'h79_79_79_79_79_79_79_79_79_79_79_79_78_78_78_78_78_78_78_78_78_78_78_78_78_78_78_77_77_77_77_77), 
	.INIT_19(256'h7C_7B_7B_7B_7B_7B_7B_7B_7B_7B_7B_7B_7B_7B_7B_7A_7A_7A_7A_7A_7A_7A_7A_7A_7A_7A_7A_7A_7A_7A_79_79), 
	.INIT_1A(256'h7E_7E_7E_7D_7D_7D_7D_7D_7D_7D_7D_7D_7D_7D_7D_7D_7D_7D_7C_7C_7C_7C_7C_7C_7C_7C_7C_7C_7C_7C_7C_7C), 
	.INIT_1B(256'h80_80_80_80_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7F_7E_7E_7E_7E_7E_7E_7E_7E_7E_7E_7E_7E), 
	.INIT_1C(256'h82_82_82_82_82_81_81_81_81_81_81_81_81_81_81_81_81_81_81_81_81_80_80_80_80_80_80_80_80_80_80_80), 
	.INIT_1D(256'h84_84_84_84_84_84_83_83_83_83_83_83_83_83_83_83_83_83_83_83_83_82_82_82_82_82_82_82_82_82_82_82), 
	.INIT_1E(256'h86_86_86_86_86_85_85_85_85_85_85_85_85_85_85_85_85_85_85_85_85_85_84_84_84_84_84_84_84_84_84_84), 
	.INIT_1F(256'h88_88_88_88_88_87_87_87_87_87_87_87_87_87_87_87_87_87_87_87_87_86_86_86_86_86_86_86_86_86_86_86), 
	// Address 1024 to 1535
	.INIT_20(256'h8A_8A_8A_89_89_89_89_89_89_89_89_89_89_89_89_89_89_89_89_89_88_88_88_88_88_88_88_88_88_88_88_88), 
	.INIT_21(256'h8C_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8B_8A_8A_8A_8A_8A_8A_8A_8A_8A_8A_8A_8A_8A_8A), 
	.INIT_22(256'h8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8D_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C_8C), 
	.INIT_23(256'h8F_8F_8F_8F_8F_8F_8F_8F_8F_8F_8F_8F_8F_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8E_8D), 
	.INIT_24(256'h91_91_91_91_91_91_91_91_91_91_90_90_90_90_90_90_90_90_90_90_90_90_90_90_90_90_90_90_8F_8F_8F_8F), 
	.INIT_25(256'h93_93_93_93_93_93_92_92_92_92_92_92_92_92_92_92_92_92_92_92_92_92_92_92_91_91_91_91_91_91_91_91), 
	.INIT_26(256'h95_94_94_94_94_94_94_94_94_94_94_94_94_94_94_94_94_94_94_93_93_93_93_93_93_93_93_93_93_93_93_93), 
	.INIT_27(256'h96_96_96_96_96_96_96_96_96_96_96_96_96_96_96_95_95_95_95_95_95_95_95_95_95_95_95_95_95_95_95_95), 
	.INIT_28(256'h98_98_98_98_98_98_98_98_98_97_97_97_97_97_97_97_97_97_97_97_97_97_97_97_97_97_97_97_96_96_96_96), 
	.INIT_29(256'h9A_9A_9A_99_99_99_99_99_99_99_99_99_99_99_99_99_99_99_99_99_99_99_98_98_98_98_98_98_98_98_98_98), 
	.INIT_2A(256'h9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9B_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A_9A), 
	.INIT_2B(256'h9D_9D_9D_9D_9D_9D_9D_9D_9D_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9C_9B_9B_9B_9B), 
	.INIT_2C(256'h9F_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9E_9D_9D_9D_9D_9D_9D_9D_9D_9D_9D_9D), 
	.INIT_2D(256'hA0_A0_A0_A0_A0_A0_A0_A0_A0_A0_A0_A0_A0_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F_9F), 
	.INIT_2E(256'hA2_A2_A2_A2_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A1_A0_A0_A0_A0_A0_A0_A0), 
	.INIT_2F(256'hA3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A3_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2_A2), 
	// Address 1536 to 2047
	.INIT_30(256'hA5_A5_A5_A5_A5_A5_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A4_A3_A3_A3_A3_A3), 
	.INIT_31(256'hA6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A6_A5_A5_A5_A5_A5_A5_A5_A5_A5_A5_A5_A5_A5_A5_A5), 
	.INIT_32(256'hA8_A8_A8_A8_A8_A8_A8_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A7_A6_A6_A6_A6), 
	.INIT_33(256'hA9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A9_A8_A8_A8_A8_A8_A8_A8_A8_A8_A8_A8_A8_A8_A8), 
	.INIT_34(256'hAB_AB_AB_AB_AB_AB_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_AA_A9_A9_A9_A9), 
	.INIT_35(256'hAC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AC_AB_AB_AB_AB_AB_AB_AB_AB_AB_AB_AB_AB_AB_AB_AB), 
	.INIT_36(256'hAE_AE_AE_AE_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AD_AC_AC_AC_AC_AC_AC), 
	.INIT_37(256'hAF_AF_AF_AF_AF_AF_AF_AF_AF_AF_AF_AF_AF_AF_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE_AE), 
	.INIT_38(256'hB1_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_B0_AF_AF_AF_AF_AF_AF_AF_AF_AF), 
	.INIT_39(256'hB2_B2_B2_B2_B2_B2_B2_B2_B2_B2_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1_B1), 
	.INIT_3A(256'hB3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B3_B2_B2_B2_B2_B2_B2_B2_B2_B2_B2_B2_B2_B2), 
	.INIT_3B(256'hB5_B5_B5_B5_B5_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B4_B3_B3_B3_B3), 
	.INIT_3C(256'hB6_B6_B6_B6_B6_B6_B6_B6_B6_B6_B6_B6_B6_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5_B5), 
	.INIT_3D(256'hB7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B7_B6_B6_B6_B6_B6_B6_B6_B6_B6_B6), 
	.INIT_3E(256'hB9_B9_B9_B9_B9_B9_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B8_B7_B7), 
	.INIT_3F(256'hBA_BA_BA_BA_BA_BA_BA_BA_BA_BA_BA_BA_BA_BA_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9_B9), 
	.SRVAL(9'h000) // Output value upon SSR assertion
	) gammalutL (
	.CLK(CLK),    // Clock
	.ADDR(DIN[10:0]),  // 11-bit Address Input
	.DO(gamma_outL), .DOP(), 
	.DI(8'h00), .DIP(1'b0), .WE(1'b0), 
	.EN(CE), .SSR(!EN || DIN[11])
	);

// Higher half of table
RAMB16_S9 #(
	// Address 2048 to 2559
	.INIT_00(256'hBB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BB_BA_BA_BA_BA_BA_BA_BA_BA_BA_BA), 
	.INIT_01(256'hBD_BD_BD_BD_BD_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BC_BB_BB), 
	.INIT_02(256'hBE_BE_BE_BE_BE_BE_BE_BE_BE_BE_BE_BE_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD_BD), 
	.INIT_03(256'hBF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BF_BE_BE_BE_BE_BE_BE_BE_BE_BE_BE_BE_BE), 
	.INIT_04(256'hC1_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_C0_BF_BF_BF_BF_BF), 
	.INIT_05(256'hC2_C2_C2_C2_C2_C2_C2_C2_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1_C1), 
	.INIT_06(256'hC3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2_C2), 
	.INIT_07(256'hC4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C4_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3_C3), 
	.INIT_08(256'hC6_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C5_C4_C4_C4_C4_C4), 
	.INIT_09(256'hC7_C7_C7_C7_C7_C7_C7_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6_C6), 
	.INIT_0A(256'hC8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7_C7), 
	.INIT_0B(256'hC9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C9_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8_C8), 
	.INIT_0C(256'hCA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_CA_C9_C9_C9_C9_C9_C9_C9_C9), 
	.INIT_0D(256'hCC_CC_CC_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CB_CA_CA_CA), 
	.INIT_0E(256'hCD_CD_CD_CD_CD_CD_CD_CD_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC_CC), 
	.INIT_0F(256'hCE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD_CD), 
	// Address 2560 to 3071
	.INIT_10(256'hCF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE_CE), 
	.INIT_11(256'hD0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_D0_CF_CF_CF_CF_CF_CF_CF_CF_CF_CF), 
	.INIT_12(256'hD1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D1_D0_D0_D0_D0_D0_D0), 
	.INIT_13(256'hD3_D3_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D2_D1_D1), 
	.INIT_14(256'hD4_D4_D4_D4_D4_D4_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3_D3), 
	.INIT_15(256'hD5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4_D4), 
	.INIT_16(256'hD6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5_D5), 
	.INIT_17(256'hD7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6_D6), 
	.INIT_18(256'hD8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D8_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7_D7), 
	.INIT_19(256'hD9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D9_D8_D8_D8_D8_D8_D8_D8_D8_D8), 
	.INIT_1A(256'hDA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_DA_D9_D9_D9_D9_D9_D9), 
	.INIT_1B(256'hDB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DB_DA_DA_DA_DA), 
	.INIT_1C(256'hDD_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DC_DB), 
	.INIT_1D(256'hDE_DE_DE_DE_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD_DD), 
	.INIT_1E(256'hDF_DF_DF_DF_DF_DF_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE_DE), 
	.INIT_1F(256'hE0_E0_E0_E0_E0_E0_E0_E0_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF_DF), 
	// Address 3072 to 3583
	.INIT_20(256'hE1_E1_E1_E1_E1_E1_E1_E1_E1_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0), 
	.INIT_21(256'hE2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1_E1), 
	.INIT_22(256'hE3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2_E2), 
	.INIT_23(256'hE4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3_E3), 
	.INIT_24(256'hE5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4_E4), 
	.INIT_25(256'hE6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5_E5), 
	.INIT_26(256'hE7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6_E6), 
	.INIT_27(256'hE8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7_E7), 
	.INIT_28(256'hE9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8_E8), 
	.INIT_29(256'hEA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9_E9), 
	.INIT_2A(256'hEB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA_EA), 
	.INIT_2B(256'hEC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB_EB), 
	.INIT_2C(256'hED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC_EC), 
	.INIT_2D(256'hEE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED_ED), 
	.INIT_2E(256'hEF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE_EE), 
	.INIT_2F(256'hF0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF_EF), 
	// Address 3584 to 4095
	.INIT_30(256'hF1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0_F0), 
	.INIT_31(256'hF2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1_F1), 
	.INIT_32(256'hF3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2_F2), 
	.INIT_33(256'hF4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3_F3), 
	.INIT_34(256'hF5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4_F4), 
	.INIT_35(256'hF6_F6_F6_F6_F6_F6_F6_F6_F6_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5_F5), 
	.INIT_36(256'hF7_F7_F7_F7_F7_F7_F7_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6_F6), 
	.INIT_37(256'hF8_F8_F8_F8_F8_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7_F7), 
	.INIT_38(256'hF9_F9_F9_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8_F8), 
	.INIT_39(256'hF9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9_F9), 
	.INIT_3A(256'hFA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA_FA), 
	.INIT_3B(256'hFB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FB_FA_FA), 
	.INIT_3C(256'hFC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FC_FB_FB_FB_FB_FB), 
	.INIT_3D(256'hFD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FC_FC_FC_FC_FC_FC_FC_FC), 
	.INIT_3E(256'hFE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD_FD), 
	.INIT_3F(256'hFF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FF_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE_FE), 
	.SRVAL(9'h000) // Output value upon SSR assertion
	) gammalutH (
	.CLK(CLK),    // Clock
	.ADDR(DIN[10:0]),  // 11-bit Address Input
	.DO(gamma_outH), .DOP(), 
	.DI(8'h00), .DIP(1'b0), .WE(1'b0), 
	.EN(CE), .SSR(!EN || !DIN[11]) // use SSR so simple OR for mux
	);

reg 	[7:0]	din_dly; // for !EN mode
always @(posedge CLK) if (CE)
	begin
	din_dly <= !EN ? DIN[11:4] : 8'h00; // make zero if enabled
	DOUT <= din_dly | gamma_outL | gamma_outH; // OR together - individually zeroed
	end


endmodule
